/*------------------------------------------------------------------------------
 Project      : IL2234 Project - Milestone 2 -> Register File 
 File         : rf_tb.sv
 Author       : Michael Kirchhofer, Yaowen Fan, Fredrik Kis
 Description  : Testbench for the processor Register File (Milestone 2).
------------------------------------------------------------------------------*/